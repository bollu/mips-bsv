module mkProc(Proc);
    Reg#(Addr) pc <- mkRegU;
